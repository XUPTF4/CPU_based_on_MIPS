module InstMem(
        input         ce,
        input  [31:0] addr,
        output  [31:0] data
    );

    reg [31:0] mem [0:1023]; // 4KB

    initial begin
        mem[0]  = 32'h0000f025;
        mem[1]  = 32'h241d1000;
        mem[2]  = 32'h8f990018;
        mem[3]  = 32'h04110038;
        mem[4]  = 32'h00000000;
        mem[5]  = 32'h00000000;
        mem[6]  = 32'h00000000;
        mem[7]  = 32'h00000000;
        mem[8]  = 32'h03a0d825;
        mem[9]  = 32'h27bdff7c;
        mem[10]  = 32'hafa10004;
        mem[11]  = 32'hafa20008;
        mem[12]  = 32'hafa3000c;
        mem[13]  = 32'hafa40010;
        mem[14]  = 32'hafa50014;
        mem[15]  = 32'hafa60018;
        mem[16]  = 32'hafa7001c;
        mem[17]  = 32'hafa80020;
        mem[18]  = 32'hafa90024;
        mem[19]  = 32'hafaa0028;
        mem[20]  = 32'hafab002c;
        mem[21]  = 32'hafac0030;
        mem[22]  = 32'hafad0034;
        mem[23]  = 32'hafae0038;
        mem[24]  = 32'hafaf003c;
        mem[25]  = 32'hafb00040;
        mem[26]  = 32'hafb10044;
        mem[27]  = 32'hafb20048;
        mem[28]  = 32'hafb3004c;
        mem[29]  = 32'hafb40050;
        mem[30]  = 32'hafb50054;
        mem[31]  = 32'hafb60058;
        mem[32]  = 32'hafb7005c;
        mem[33]  = 32'hafb80060;
        mem[34]  = 32'hafb90064;
        mem[35]  = 32'hafbc0070;
        mem[36]  = 32'hafbe0078;
        mem[37]  = 32'hafbf007c;
        mem[38]  = 32'hafbb0074;
        mem[39]  = 32'h03a02025;
        mem[40]  = 32'h8f99001c;
        mem[41]  = 32'h0411003c;
        mem[42]  = 32'h00000000;
        mem[43]  = 32'h8c440010;
        mem[44]  = 32'h8c480080;
        mem[45]  = 32'h00000000;
        mem[46]  = 32'h00000000;
        mem[47]  = 32'h00000000;
        mem[48]  = 32'h00000000;
        mem[49]  = 32'h00000000;
        mem[50]  = 32'h40880000;
        mem[51]  = 32'h27bd0084;
        mem[52]  = 32'h42000018;
        mem[53]  = 32'h00000000;
        mem[54]  = 32'h00000000;
        mem[55]  = 32'h00000000;
        mem[56]  = 32'h00802025;
        mem[57]  = 32'h0000000d;
        mem[58]  = 32'h1000ffff;
        mem[59]  = 32'h00000000;
        mem[60]  = 32'h3c1c0000;
        mem[61]  = 32'h279c0000;
        mem[62]  = 32'h27bdffe0;
        mem[63]  = 32'h8f990020;
        mem[64]  = 32'hafbf001c;
        mem[65]  = 32'hafbc0010;
        mem[66]  = 32'h04110045;
        mem[67]  = 32'h00000000;
        mem[68]  = 32'h00402025;
        mem[69]  = 32'h0c000038;
        mem[70]  = 32'h00000000;
        mem[71]  = 32'h00000000;
        mem[72]  = 32'h10800003;
        mem[73]  = 32'h00000000;
        mem[74]  = 32'h03e00008;
        mem[75]  = 32'h00000000;
        mem[76]  = 32'h3c1c0000;
        mem[77]  = 32'h279c0000;
        mem[78]  = 32'h8f990024;
        mem[79]  = 32'h24040001;
        mem[80]  = 32'h1000ffe7;
        mem[81]  = 32'h00000000;
        mem[82]  = 32'h0000000c;
        mem[83]  = 32'h00000000;
        mem[84]  = 32'h03e00008;
        mem[85]  = 32'h00000000;
        mem[86]  = 32'h3c030000;
        mem[87]  = 32'h8c620030;
        mem[88]  = 32'h00000000;
        mem[89]  = 32'h24420001;
        mem[90]  = 32'h30440001;
        mem[91]  = 32'hac620030;
        mem[92]  = 32'h14800005;
        mem[93]  = 32'h00000000;
        mem[94]  = 32'h3c020000;
        mem[95]  = 32'h8c4200b8;
        mem[96]  = 32'h03e00008;
        mem[97]  = 32'h00000000;
        mem[98]  = 32'h3c020000;
        mem[99]  = 32'h8c42013c;
        mem[100]  = 32'h03e00008;
        mem[101]  = 32'h00000000;
        mem[102]  = 32'h08000056;
        mem[103]  = 32'h00000000;
        mem[104]  = 32'hafa40000;
        mem[105]  = 32'hafa50004;
        mem[106]  = 32'haca7ff8c;
        mem[107]  = 32'haca6fffc;
        mem[108]  = 32'h24a2ff7c;
        mem[109]  = 32'h03e00008;
        mem[110]  = 32'h00000000;
        mem[111]  = 32'hac040ffc;
        mem[112]  = 32'hac040ff8;
        mem[113]  = 32'h03e00008;
        mem[114]  = 32'h00000000;
        mem[115]  = 32'h27bdffe0;
        mem[116]  = 32'h3c065555;
        mem[117]  = 32'h3c02aaaa;
        mem[118]  = 32'h00801825;
        mem[119]  = 32'hafbf001c;
        mem[120]  = 32'h24050001;
        mem[121]  = 32'h24c65555;
        mem[122]  = 32'h3442aaaa;
        mem[123]  = 32'h00402025;
        mem[124]  = 32'h10650002;
        mem[125]  = 32'h00000000;
        mem[126]  = 32'h00c02025;
        mem[127]  = 32'h0c00006f;
        mem[128]  = 32'h00000000;
        mem[129]  = 32'h0c000052;
        mem[130]  = 32'h00000000;
        mem[131]  = 32'h1000fff7;
        mem[132]  = 32'h00000000;
        mem[133]  = 32'h00000000;
        mem[134]  = 32'h00000000;
        mem[135]  = 32'h00000000;
        mem[136]  = 32'h3c080000;
        mem[137]  = 32'h250300b8;
        mem[138]  = 32'h3c050000;
        mem[139]  = 32'h3c060000;
        mem[140]  = 32'h27bdffd0;
        mem[141]  = 32'h24c601cc;
        mem[142]  = 32'h00602025;
        mem[143]  = 32'h24a5013c;
        mem[144]  = 32'h24070001;
        mem[145]  = 32'hafbf002c;
        mem[146]  = 32'h0c000068;
        mem[147]  = 32'h00000000;
        mem[148]  = 32'h00a02025;
        mem[149]  = 32'h3c050000;
        mem[150]  = 32'h24070002;
        mem[151]  = 32'h24a501c0;
        mem[152]  = 32'had0200b8;
        mem[153]  = 32'h0c000068;
        mem[154]  = 32'h00000000;
        mem[155]  = 32'hac620084;
        mem[156]  = 32'h00002025;
        mem[157]  = 32'h0c000052;
        mem[158]  = 32'h00000000;
        mem[159]  = 32'h0c000048;
        mem[160]  = 32'h00000000;
        mem[161]  = 32'h8fbf002c;
        mem[162]  = 32'h00001025;
        mem[163]  = 32'h27bd0030;
        mem[164]  = 32'h03e00008;
        mem[165]  = 32'h00000000;
    end
    assign data = ce ? mem[addr >> 2] : 32'b0;

endmodule
