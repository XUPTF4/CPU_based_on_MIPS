module InstMem(
        input         ce,
        input  [31:0] addr,
        output  [31:0] data
    );

    reg [31:0] mem [0:1023]; // 4KB

    initial begin
        mem[0]  = 32'h0000f025;
        mem[1]  = 32'h241d1000;
        mem[2]  = 32'h8f990148;
        mem[3]  = 32'h04110038;
        mem[4]  = 32'h00000000;
        mem[5]  = 32'h00000000;
        mem[6]  = 32'h00000000;
        mem[7]  = 32'h00000000;
        mem[8]  = 32'h10800003;
        mem[9]  = 32'h00000000;
        mem[10]  = 32'h03e00008;
        mem[11]  = 32'h00000000;
        mem[12]  = 32'h3c1c0000;
        mem[13]  = 32'h279c0000;
        mem[14]  = 32'h8f99014c;
        mem[15]  = 32'h24040001;
        mem[16]  = 32'h10000027;
        mem[17]  = 32'h00000000;
        mem[18]  = 32'h00000000;
        mem[19]  = 32'h00000000;
        mem[20]  = 32'h27bdffd8;
        mem[21]  = 32'hafb00018;
        mem[22]  = 32'h3c100000;
        mem[23]  = 32'hafb1001c;
        mem[24]  = 32'h261000a0;
        mem[25]  = 32'h3c110000;
        mem[26]  = 32'hafb20020;
        mem[27]  = 32'hafbf0024;
        mem[28]  = 32'h26310008;
        mem[29]  = 32'h26120098;
        mem[30]  = 32'h8e020004;
        mem[31]  = 32'h8e030000;
        mem[32]  = 32'h8e240000;
        mem[33]  = 32'h00431021;
        mem[34]  = 32'h00822026;
        mem[35]  = 32'hae020008;
        mem[36]  = 32'h2c840001;
        mem[37]  = 32'h26100004;
        mem[38]  = 32'h0c000008;
        mem[39]  = 32'h00000000;
        mem[40]  = 32'h26310004;
        mem[41]  = 32'h1612fff4;
        mem[42]  = 32'h00000000;
        mem[43]  = 32'h24040001;
        mem[44]  = 32'h0c000008;
        mem[45]  = 32'h00000000;
        mem[46]  = 32'h8fbf0024;
        mem[47]  = 32'h8fb20020;
        mem[48]  = 32'h8fb1001c;
        mem[49]  = 32'h8fb00018;
        mem[50]  = 32'h00001025;
        mem[51]  = 32'h27bd0028;
        mem[52]  = 32'h03e00008;
        mem[53]  = 32'h00000000;
        mem[54]  = 32'h00000000;
        mem[55]  = 32'h00000000;
        mem[56]  = 32'h00802025;
        mem[57]  = 32'h0000000d;
        mem[58]  = 32'h1000ffff;
        mem[59]  = 32'h00000000;
        mem[60]  = 32'h3c1c0000;
        mem[61]  = 32'h279c0000;
        mem[62]  = 32'h27bdffe0;
        mem[63]  = 32'h8f990150;
        mem[64]  = 32'hafbf001c;
        mem[65]  = 32'hafbc0010;
        mem[66]  = 32'h0411ffd1;
        mem[67]  = 32'h00000000;
        mem[68]  = 32'h00402025;
        mem[69]  = 32'h0000000d;
        mem[70]  = 32'h1000ffff;
        mem[71]  = 32'h00000000;
    end
    assign data = ce ? mem[addr >> 2] : 32'b0;

endmodule
