module InstMem(
        input         ce,
        input  [31:0] addr,
        output  [31:0] data
    );

    reg [31:0] mem [0:1023]; // 4KB

    initial begin
        mem[0]  = 32'h0000f025;
        mem[1]  = 32'h241d1000;
        mem[2]  = 32'h8f990038;
        mem[3]  = 32'h04110044;
        mem[4]  = 32'h00000000;
        mem[5]  = 32'h00000000;
        mem[6]  = 32'h00000000;
        mem[7]  = 32'h00000000;
        mem[8]  = 32'h10800003;
        mem[9]  = 32'h00000000;
        mem[10]  = 32'h03e00008;
        mem[11]  = 32'h00000000;
        mem[12]  = 32'h3c1c0000;
        mem[13]  = 32'h279c0000;
        mem[14]  = 32'h8f99003c;
        mem[15]  = 32'h24040001;
        mem[16]  = 32'h10000033;
        mem[17]  = 32'h00000000;
        mem[18]  = 32'h00000000;
        mem[19]  = 32'h00000000;
        mem[20]  = 32'h27bdffd0;
        mem[21]  = 32'hafb10020;
        mem[22]  = 32'h3c110000;
        mem[23]  = 32'hafb30028;
        mem[24]  = 32'hafb20024;
        mem[25]  = 32'hafb0001c;
        mem[26]  = 32'hafbf002c;
        mem[27]  = 32'h00009025;
        mem[28]  = 32'h24100065;
        mem[29]  = 32'h26310000;
        mem[30]  = 32'h24130097;
        mem[31]  = 32'h24020002;
        mem[32]  = 32'h0202001a;
        mem[33]  = 32'h14400002;
        mem[34]  = 32'h00000000;
        mem[35]  = 32'h0007000d;
        mem[36]  = 32'h24420001;
        mem[37]  = 32'h00001810;
        mem[38]  = 32'h1060000b;
        mem[39]  = 32'h00000000;
        mem[40]  = 32'h1450fff7;
        mem[41]  = 32'h00000000;
        mem[42]  = 32'h00121080;
        mem[43]  = 32'h00511021;
        mem[44]  = 32'h8c440000;
        mem[45]  = 32'h26520001;
        mem[46]  = 32'h00902026;
        mem[47]  = 32'h2c840001;
        mem[48]  = 32'h0c000008;
        mem[49]  = 32'h00000000;
        mem[50]  = 32'h26100002;
        mem[51]  = 32'h1613ffeb;
        mem[52]  = 32'h00000000;
        mem[53]  = 32'h3a44000a;
        mem[54]  = 32'h2c840001;
        mem[55]  = 32'h0c000008;
        mem[56]  = 32'h00000000;
        mem[57]  = 32'h8fbf002c;
        mem[58]  = 32'h8fb30028;
        mem[59]  = 32'h8fb20024;
        mem[60]  = 32'h8fb10020;
        mem[61]  = 32'h8fb0001c;
        mem[62]  = 32'h00001025;
        mem[63]  = 32'h27bd0030;
        mem[64]  = 32'h03e00008;
        mem[65]  = 32'h00000000;
        mem[66]  = 32'h00000000;
        mem[67]  = 32'h00000000;
        mem[68]  = 32'h00802025;
        mem[69]  = 32'h0000000d;
        mem[70]  = 32'h1000ffff;
        mem[71]  = 32'h00000000;
        mem[72]  = 32'h3c1c0000;
        mem[73]  = 32'h279c0000;
        mem[74]  = 32'h27bdffe0;
        mem[75]  = 32'h8f990040;
        mem[76]  = 32'hafbf001c;
        mem[77]  = 32'hafbc0010;
        mem[78]  = 32'h0411ffc5;
        mem[79]  = 32'h00000000;
        mem[80]  = 32'h00402025;
        mem[81]  = 32'h0000000d;
        mem[82]  = 32'h1000ffff;
        mem[83]  = 32'h00000000;
    end
    assign data = ce ? mem[addr >> 2] : 32'b0;

endmodule
