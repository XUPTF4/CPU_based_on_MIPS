module InstMem(
        input         ce,
        input  [31:0] addr,
        output  [31:0] data
    );

    reg [31:0] mem [0:1023]; // 4KB

    initial begin
        mem[0]  = 32'h0000f025;
        mem[1]  = 32'h241d1000;
        mem[2]  = 32'h8f990008;
        mem[3]  = 32'h04110086;
        mem[4]  = 32'h00000000;
        mem[5]  = 32'h00000000;
        mem[6]  = 32'h00000000;
        mem[7]  = 32'h00000000;
        mem[8]  = 32'h27bdffe0;
        mem[9]  = 32'hafbf001c;
        mem[10]  = 32'hafbe0018;
        mem[11]  = 32'h03a0f025;
        mem[12]  = 32'h3c1c0000;
        mem[13]  = 32'h279c0000;
        mem[14]  = 32'hafbc0010;
        mem[15]  = 32'hafc40020;
        mem[16]  = 32'h8fc20020;
        mem[17]  = 32'h00000000;
        mem[18]  = 32'h14400008;
        mem[19]  = 32'h00000000;
        mem[20]  = 32'h24040001;
        mem[21]  = 32'h8f82000c;
        mem[22]  = 32'h00000000;
        mem[23]  = 32'h0040c825;
        mem[24]  = 32'h04110067;
        mem[25]  = 32'h00000000;
        mem[26]  = 32'h8fdc0010;
        mem[27]  = 32'h00000000;
        mem[28]  = 32'h03c0e825;
        mem[29]  = 32'h8fbf001c;
        mem[30]  = 32'h8fbe0018;
        mem[31]  = 32'h27bd0020;
        mem[32]  = 32'h03e00008;
        mem[33]  = 32'h00000000;
        mem[34]  = 32'h27bdffd0;
        mem[35]  = 32'hafbf002c;
        mem[36]  = 32'hafbe0028;
        mem[37]  = 32'h03a0f025;
        mem[38]  = 32'h2402000a;
        mem[39]  = 32'hafc2001c;
        mem[40]  = 32'h24020005;
        mem[41]  = 32'hafc20020;
        mem[42]  = 32'h8fc3001c;
        mem[43]  = 32'h8fc20020;
        mem[44]  = 32'h00000000;
        mem[45]  = 32'h00621021;
        mem[46]  = 32'hafc20024;
        mem[47]  = 32'h8fc20024;
        mem[48]  = 32'h00000000;
        mem[49]  = 32'h3842000f;
        mem[50]  = 32'h2c420001;
        mem[51]  = 32'h304200ff;
        mem[52]  = 32'h00402025;
        mem[53]  = 32'h0c000008;
        mem[54]  = 32'h00000000;
        mem[55]  = 32'h8fc3001c;
        mem[56]  = 32'h8fc20020;
        mem[57]  = 32'h00000000;
        mem[58]  = 32'h00621023;
        mem[59]  = 32'hafc20024;
        mem[60]  = 32'h8fc20024;
        mem[61]  = 32'h00000000;
        mem[62]  = 32'h38420005;
        mem[63]  = 32'h2c420001;
        mem[64]  = 32'h304200ff;
        mem[65]  = 32'h00402025;
        mem[66]  = 32'h0c000008;
        mem[67]  = 32'h00000000;
        mem[68]  = 32'h8fc20024;
        mem[69]  = 32'h00000000;
        mem[70]  = 32'h1840000a;
        mem[71]  = 32'h00000000;
        mem[72]  = 32'h8fc20024;
        mem[73]  = 32'h00000000;
        mem[74]  = 32'h0002102a;
        mem[75]  = 32'h304200ff;
        mem[76]  = 32'h00402025;
        mem[77]  = 32'h0c000008;
        mem[78]  = 32'h00000000;
        mem[79]  = 32'h10000015;
        mem[80]  = 32'h00000000;
        mem[81]  = 32'h8fc20024;
        mem[82]  = 32'h00000000;
        mem[83]  = 32'h0441000a;
        mem[84]  = 32'h00000000;
        mem[85]  = 32'h8fc20024;
        mem[86]  = 32'h00000000;
        mem[87]  = 32'h000217c2;
        mem[88]  = 32'h304200ff;
        mem[89]  = 32'h00402025;
        mem[90]  = 32'h0c000008;
        mem[91]  = 32'h00000000;
        mem[92]  = 32'h10000008;
        mem[93]  = 32'h00000000;
        mem[94]  = 32'h8fc20024;
        mem[95]  = 32'h00000000;
        mem[96]  = 32'h2c420001;
        mem[97]  = 32'h304200ff;
        mem[98]  = 32'h00402025;
        mem[99]  = 32'h0c000008;
        mem[100]  = 32'h00000000;
        mem[101]  = 32'hafc00018;
        mem[102]  = 32'h10000005;
        mem[103]  = 32'h00000000;
        mem[104]  = 32'h8fc20018;
        mem[105]  = 32'h00000000;
        mem[106]  = 32'h24420001;
        mem[107]  = 32'hafc20018;
        mem[108]  = 32'h8fc20018;
        mem[109]  = 32'h00000000;
        mem[110]  = 32'h28420005;
        mem[111]  = 32'h1440fff8;
        mem[112]  = 32'h00000000;
        mem[113]  = 32'h8fc20018;
        mem[114]  = 32'h00000000;
        mem[115]  = 32'h38420005;
        mem[116]  = 32'h2c420001;
        mem[117]  = 32'h304200ff;
        mem[118]  = 32'h00402025;
        mem[119]  = 32'h0c000008;
        mem[120]  = 32'h00000000;
        mem[121]  = 32'h00001025;
        mem[122]  = 32'h03c0e825;
        mem[123]  = 32'h8fbf002c;
        mem[124]  = 32'h8fbe0028;
        mem[125]  = 32'h27bd0030;
        mem[126]  = 32'h03e00008;
        mem[127]  = 32'h00000000;
        mem[128]  = 32'h27bdfff8;
        mem[129]  = 32'hafbe0004;
        mem[130]  = 32'h03a0f025;
        mem[131]  = 32'hafc40008;
        mem[132]  = 32'h8fc20008;
        mem[133]  = 32'h00000000;
        mem[134]  = 32'h00402025;
        mem[135]  = 32'h0000000d;
        mem[136]  = 32'h1000ffff;
        mem[137]  = 32'h00000000;
        mem[138]  = 32'h27bdffd8;
        mem[139]  = 32'hafbf0024;
        mem[140]  = 32'hafbe0020;
        mem[141]  = 32'h03a0f025;
        mem[142]  = 32'h3c1c0000;
        mem[143]  = 32'h279c0000;
        mem[144]  = 32'hafbc0010;
        mem[145]  = 32'h8f820010;
        mem[146]  = 32'h00000000;
        mem[147]  = 32'h0040c825;
        mem[148]  = 32'h0411ff8d;
        mem[149]  = 32'h00000000;
        mem[150]  = 32'h8fdc0010;
        mem[151]  = 32'hafc20018;
        mem[152]  = 32'h8fc40018;
        mem[153]  = 32'h0c000080;
        mem[154]  = 32'h00000000;
        mem[155]  = 32'h8fdc0010;
        mem[156]  = 32'h00000000;
        mem[157]  = 32'h03c0e825;
        mem[158]  = 32'h8fbf0024;
        mem[159]  = 32'h8fbe0020;
        mem[160]  = 32'h27bd0028;
        mem[161]  = 32'h03e00008;
        mem[162]  = 32'h00000000;
        mem[163]  = 32'h00000000;
    end
    assign data = ce ? mem[addr >> 2] : 32'b0;

endmodule
