module InstMem(
        input         ce,
        input  [31:0] addr,
        output  [31:0] data
    );

    reg [31:0] mem [0:1023]; // 4KB

    initial begin
        mem[0]  = 32'h0000f025;
        mem[1]  = 32'h241d1000;
        mem[2]  = 32'h8f990068;
        mem[3]  = 32'h04110060;
        mem[4]  = 32'h00000000;
        mem[5]  = 32'h00000000;
        mem[6]  = 32'h00000000;
        mem[7]  = 32'h00000000;
        mem[8]  = 32'h10800003;
        mem[9]  = 32'h00000000;
        mem[10]  = 32'h03e00008;
        mem[11]  = 32'h00000000;
        mem[12]  = 32'h3c1c0000;
        mem[13]  = 32'h279c0000;
        mem[14]  = 32'h8f99006c;
        mem[15]  = 32'h24040001;
        mem[16]  = 32'h1000004f;
        mem[17]  = 32'h00000000;
        mem[18]  = 32'h00870018;
        mem[19]  = 32'h00002012;
        mem[20]  = 32'h00000000;
        mem[21]  = 32'h00000000;
        mem[22]  = 32'h00c50018;
        mem[23]  = 32'h00003012;
        mem[24]  = 32'h00862021;
        mem[25]  = 32'h00000000;
        mem[26]  = 32'h00a70019;
        mem[27]  = 32'h00001010;
        mem[28]  = 32'h00821021;
        mem[29]  = 32'h00001812;
        mem[30]  = 32'h03e00008;
        mem[31]  = 32'h00000000;
        mem[32]  = 32'h27bdffc0;
        mem[33]  = 32'hafb70038;
        mem[34]  = 32'hafb4002c;
        mem[35]  = 32'h3c170000;
        mem[36]  = 32'h3c140000;
        mem[37]  = 32'hafb30028;
        mem[38]  = 32'hafb20024;
        mem[39]  = 32'hafb10020;
        mem[40]  = 32'hafbf003c;
        mem[41]  = 32'hafb60034;
        mem[42]  = 32'hafb50030;
        mem[43]  = 32'hafb0001c;
        mem[44]  = 32'h26f70050;
        mem[45]  = 32'h00009025;
        mem[46]  = 32'h00008825;
        mem[47]  = 32'h26940000;
        mem[48]  = 32'h24130004;
        mem[49]  = 32'h001280c0;
        mem[50]  = 32'h02908021;
        mem[51]  = 32'h02e0b025;
        mem[52]  = 32'h0220a825;
        mem[53]  = 32'h8ec20000;
        mem[54]  = 32'h8ee30000;
        mem[55]  = 32'h8e040000;
        mem[56]  = 32'h00620018;
        mem[57]  = 32'h8e020004;
        mem[58]  = 32'h26b50001;
        mem[59]  = 32'h26100008;
        mem[60]  = 32'h26d60004;
        mem[61]  = 32'h00003812;
        mem[62]  = 32'h00471026;
        mem[63]  = 32'h00003010;
        mem[64]  = 32'h00862026;
        mem[65]  = 32'h00822025;
        mem[66]  = 32'h2c840001;
        mem[67]  = 32'h0c000008;
        mem[68]  = 32'h00000000;
        mem[69]  = 32'h16b3ffef;
        mem[70]  = 32'h00000000;
        mem[71]  = 32'h26520004;
        mem[72]  = 32'h02519023;
        mem[73]  = 32'h24040001;
        mem[74]  = 32'h26310001;
        mem[75]  = 32'h0c000008;
        mem[76]  = 32'h00000000;
        mem[77]  = 32'h26f70004;
        mem[78]  = 32'h1635ffe2;
        mem[79]  = 32'h00000000;
        mem[80]  = 32'h24040001;
        mem[81]  = 32'h0c000008;
        mem[82]  = 32'h00000000;
        mem[83]  = 32'h8fbf003c;
        mem[84]  = 32'h8fb70038;
        mem[85]  = 32'h8fb60034;
        mem[86]  = 32'h8fb50030;
        mem[87]  = 32'h8fb4002c;
        mem[88]  = 32'h8fb30028;
        mem[89]  = 32'h8fb20024;
        mem[90]  = 32'h8fb10020;
        mem[91]  = 32'h8fb0001c;
        mem[92]  = 32'h00001025;
        mem[93]  = 32'h27bd0040;
        mem[94]  = 32'h03e00008;
        mem[95]  = 32'h00000000;
        mem[96]  = 32'h00802025;
        mem[97]  = 32'h0000000d;
        mem[98]  = 32'h1000ffff;
        mem[99]  = 32'h00000000;
        mem[100]  = 32'h3c1c0000;
        mem[101]  = 32'h279c0000;
        mem[102]  = 32'h27bdffe0;
        mem[103]  = 32'h8f990070;
        mem[104]  = 32'hafbf001c;
        mem[105]  = 32'hafbc0010;
        mem[106]  = 32'h0411ffb5;
        mem[107]  = 32'h00000000;
        mem[108]  = 32'h00402025;
        mem[109]  = 32'h0000000d;
        mem[110]  = 32'h1000ffff;
        mem[111]  = 32'h00000000;
    end
    assign data = ce ? mem[addr >> 2] : 32'b0;

endmodule
