module InstMem(
        input         ce,
        input  [31:0] addr,
        output  [31:0] data
    );

    reg [31:0] mem [0:1023]; // 4KB

    initial begin
        mem[0]  = 32'h0000f025;
        mem[1]  = 32'h241d1000;
        mem[2]  = 32'h8f990018;
        mem[3]  = 32'h0411003e;
        mem[4]  = 32'h00000000;
        mem[5]  = 32'h00000000;
        mem[6]  = 32'h00000000;
        mem[7]  = 32'h00000000;
        mem[8]  = 32'h03a0d825;
        mem[9]  = 32'h27bdff7c;
        mem[10]  = 32'hafa10004;
        mem[11]  = 32'hafa20008;
        mem[12]  = 32'hafa3000c;
        mem[13]  = 32'hafa40010;
        mem[14]  = 32'hafa50014;
        mem[15]  = 32'hafa60018;
        mem[16]  = 32'hafa7001c;
        mem[17]  = 32'hafa80020;
        mem[18]  = 32'hafa90024;
        mem[19]  = 32'hafaa0028;
        mem[20]  = 32'hafab002c;
        mem[21]  = 32'hafac0030;
        mem[22]  = 32'hafad0034;
        mem[23]  = 32'hafae0038;
        mem[24]  = 32'hafaf003c;
        mem[25]  = 32'hafb00040;
        mem[26]  = 32'hafb10044;
        mem[27]  = 32'hafb20048;
        mem[28]  = 32'hafb3004c;
        mem[29]  = 32'hafb40050;
        mem[30]  = 32'hafb50054;
        mem[31]  = 32'hafb60058;
        mem[32]  = 32'hafb7005c;
        mem[33]  = 32'hafb80060;
        mem[34]  = 32'hafb90064;
        mem[35]  = 32'hafbc0070;
        mem[36]  = 32'hafbe0078;
        mem[37]  = 32'hafbf007c;
        mem[38]  = 32'hafbb0074;
        mem[39]  = 32'h03a02025;
        mem[40]  = 32'h8f99001c;
        mem[41]  = 32'h04110078;
        mem[42]  = 32'h00000000;
        mem[43]  = 32'h8c440010;
        mem[44]  = 32'h8c480080;
        mem[45]  = 32'h00000000;
        mem[46]  = 32'h00000000;
        mem[47]  = 32'h00000000;
        mem[48]  = 32'h00000000;
        mem[49]  = 32'h00000000;
        mem[50]  = 32'h40880000;
        mem[51]  = 32'h27bd0084;
        mem[52]  = 32'h42000018;
        mem[53]  = 32'h00000000;
        mem[54]  = 32'h00000000;
        mem[55]  = 32'h00000000;
        mem[56]  = 32'h27bdfff8;
        mem[57]  = 32'hafbe0004;
        mem[58]  = 32'h03a0f025;
        mem[59]  = 32'hafc40008;
        mem[60]  = 32'h8fc20008;
        mem[61]  = 32'h00000000;
        mem[62]  = 32'h00402025;
        mem[63]  = 32'h0000000d;
        mem[64]  = 32'h1000ffff;
        mem[65]  = 32'h00000000;
        mem[66]  = 32'h27bdffd8;
        mem[67]  = 32'hafbf0024;
        mem[68]  = 32'hafbe0020;
        mem[69]  = 32'h03a0f025;
        mem[70]  = 32'h3c1c0000;
        mem[71]  = 32'h279c0000;
        mem[72]  = 32'hafbc0010;
        mem[73]  = 32'h8f820020;
        mem[74]  = 32'h00000000;
        mem[75]  = 32'h0040c825;
        mem[76]  = 32'h041100ab;
        mem[77]  = 32'h00000000;
        mem[78]  = 32'h8fdc0010;
        mem[79]  = 32'hafc20018;
        mem[80]  = 32'h8fc40018;
        mem[81]  = 32'h0c000038;
        mem[82]  = 32'h00000000;
        mem[83]  = 32'h8fdc0010;
        mem[84]  = 32'h00000000;
        mem[85]  = 32'h03c0e825;
        mem[86]  = 32'h8fbf0024;
        mem[87]  = 32'h8fbe0020;
        mem[88]  = 32'h27bd0028;
        mem[89]  = 32'h03e00008;
        mem[90]  = 32'h00000000;
        mem[91]  = 32'h00000000;
        mem[92]  = 32'h27bdffe0;
        mem[93]  = 32'hafbf001c;
        mem[94]  = 32'hafbe0018;
        mem[95]  = 32'h03a0f025;
        mem[96]  = 32'h3c1c0000;
        mem[97]  = 32'h279c0000;
        mem[98]  = 32'hafbc0010;
        mem[99]  = 32'hafc40020;
        mem[100]  = 32'h8fc20020;
        mem[101]  = 32'h00000000;
        mem[102]  = 32'h14400008;
        mem[103]  = 32'h00000000;
        mem[104]  = 32'h24040001;
        mem[105]  = 32'h8f820024;
        mem[106]  = 32'h00000000;
        mem[107]  = 32'h0040c825;
        mem[108]  = 32'h0411ffcb;
        mem[109]  = 32'h00000000;
        mem[110]  = 32'h8fdc0010;
        mem[111]  = 32'h00000000;
        mem[112]  = 32'h03c0e825;
        mem[113]  = 32'h8fbf001c;
        mem[114]  = 32'h8fbe0018;
        mem[115]  = 32'h27bd0020;
        mem[116]  = 32'h03e00008;
        mem[117]  = 32'h00000000;
        mem[118]  = 32'h27bdfff8;
        mem[119]  = 32'hafbe0004;
        mem[120]  = 32'h03a0f025;
        mem[121]  = 32'h0000000c;
        mem[122]  = 32'h00000000;
        mem[123]  = 32'h00000000;
        mem[124]  = 32'h03c0e825;
        mem[125]  = 32'h8fbe0004;
        mem[126]  = 32'h27bd0008;
        mem[127]  = 32'h03e00008;
        mem[128]  = 32'h00000000;
        mem[129]  = 32'h27bdffe8;
        mem[130]  = 32'hafbe0014;
        mem[131]  = 32'h03a0f025;
        mem[132]  = 32'hafc40018;
        mem[133]  = 32'h3c020000;
        mem[134]  = 32'h8c4201bc;
        mem[135]  = 32'h00000000;
        mem[136]  = 32'h24430001;
        mem[137]  = 32'h3c020000;
        mem[138]  = 32'hac4301bc;
        mem[139]  = 32'h3c020000;
        mem[140]  = 32'h8c4201bc;
        mem[141]  = 32'h00000000;
        mem[142]  = 32'h30420001;
        mem[143]  = 32'h14400007;
        mem[144]  = 32'h00000000;
        mem[145]  = 32'h3c020000;
        mem[146]  = 32'h8c420030;
        mem[147]  = 32'h00000000;
        mem[148]  = 32'hafc20008;
        mem[149]  = 32'h10000006;
        mem[150]  = 32'h00000000;
        mem[151]  = 32'h3c020000;
        mem[152]  = 32'h24420030;
        mem[153]  = 32'h8c420084;
        mem[154]  = 32'h00000000;
        mem[155]  = 32'hafc20008;
        mem[156]  = 32'h8fc20008;
        mem[157]  = 32'h03c0e825;
        mem[158]  = 32'h8fbe0014;
        mem[159]  = 32'h27bd0018;
        mem[160]  = 32'h03e00008;
        mem[161]  = 32'h00000000;
        mem[162]  = 32'h27bdffe0;
        mem[163]  = 32'hafbf001c;
        mem[164]  = 32'hafbe0018;
        mem[165]  = 32'h03a0f025;
        mem[166]  = 32'hafc40020;
        mem[167]  = 32'h8fc40020;
        mem[168]  = 32'h0c000081;
        mem[169]  = 32'h00000000;
        mem[170]  = 32'hafc20020;
        mem[171]  = 32'h8fc20020;
        mem[172]  = 32'h03c0e825;
        mem[173]  = 32'h8fbf001c;
        mem[174]  = 32'h8fbe0018;
        mem[175]  = 32'h27bd0020;
        mem[176]  = 32'h03e00008;
        mem[177]  = 32'h00000000;
        mem[178]  = 32'h27bdffe8;
        mem[179]  = 32'hafbe0014;
        mem[180]  = 32'h03a0f025;
        mem[181]  = 32'hafc40018;
        mem[182]  = 32'hafc5001c;
        mem[183]  = 32'hafc60020;
        mem[184]  = 32'hafc70024;
        mem[185]  = 32'h8fc2001c;
        mem[186]  = 32'h00000000;
        mem[187]  = 32'h2442ff7c;
        mem[188]  = 32'hafc20008;
        mem[189]  = 32'h8fc30024;
        mem[190]  = 32'h8fc20008;
        mem[191]  = 32'h00000000;
        mem[192]  = 32'hac430010;
        mem[193]  = 32'h8fc30020;
        mem[194]  = 32'h8fc20008;
        mem[195]  = 32'h00000000;
        mem[196]  = 32'hac430080;
        mem[197]  = 32'h8fc20008;
        mem[198]  = 32'h03c0e825;
        mem[199]  = 32'h8fbe0014;
        mem[200]  = 32'h27bd0018;
        mem[201]  = 32'h03e00008;
        mem[202]  = 32'h00000000;
        mem[203]  = 32'h27bdffe8;
        mem[204]  = 32'hafbe0014;
        mem[205]  = 32'h03a0f025;
        mem[206]  = 32'hafc40018;
        mem[207]  = 32'h24020ffc;
        mem[208]  = 32'hafc20008;
        mem[209]  = 32'h8fc20008;
        mem[210]  = 32'h8fc30018;
        mem[211]  = 32'h00000000;
        mem[212]  = 32'hac430000;
        mem[213]  = 32'h24020ff8;
        mem[214]  = 32'hafc2000c;
        mem[215]  = 32'h8fc2000c;
        mem[216]  = 32'h8fc30018;
        mem[217]  = 32'h00000000;
        mem[218]  = 32'hac430000;
        mem[219]  = 32'h00000000;
        mem[220]  = 32'h03c0e825;
        mem[221]  = 32'h8fbe0014;
        mem[222]  = 32'h27bd0018;
        mem[223]  = 32'h03e00008;
        mem[224]  = 32'h00000000;
        mem[225]  = 32'h27bdffe0;
        mem[226]  = 32'hafbf001c;
        mem[227]  = 32'hafbe0018;
        mem[228]  = 32'h03a0f025;
        mem[229]  = 32'hafc40020;
        mem[230]  = 32'h8fc30020;
        mem[231]  = 32'h24020001;
        mem[232]  = 32'h14620007;
        mem[233]  = 32'h00000000;
        mem[234]  = 32'h3c02aaaa;
        mem[235]  = 32'h3444aaaa;
        mem[236]  = 32'h0c0000cb;
        mem[237]  = 32'h00000000;
        mem[238]  = 32'h10000005;
        mem[239]  = 32'h00000000;
        mem[240]  = 32'h3c025555;
        mem[241]  = 32'h34445555;
        mem[242]  = 32'h0c0000cb;
        mem[243]  = 32'h00000000;
        mem[244]  = 32'h0c000076;
        mem[245]  = 32'h00000000;
        mem[246]  = 32'h1000ffef;
        mem[247]  = 32'h00000000;
        mem[248]  = 32'h27bdffd0;
        mem[249]  = 32'hafbf002c;
        mem[250]  = 32'hafbe0028;
        mem[251]  = 32'h03a0f025;
        mem[252]  = 32'h3c020000;
        mem[253]  = 32'h24420030;
        mem[254]  = 32'hafc20018;
        mem[255]  = 32'h3c020000;
        mem[256]  = 32'h244200b4;
        mem[257]  = 32'hafc2001c;
        mem[258]  = 32'h24070001;
        mem[259]  = 32'h3c020000;
        mem[260]  = 32'h24460384;
        mem[261]  = 32'h8fc40018;
        mem[262]  = 32'h8fc5001c;
        mem[263]  = 32'h0c0000b2;
        mem[264]  = 32'h00000000;
        mem[265]  = 32'h00401825;
        mem[266]  = 32'h3c020000;
        mem[267]  = 32'hac430030;
        mem[268]  = 32'h3c020000;
        mem[269]  = 32'h244200b4;
        mem[270]  = 32'hafc20020;
        mem[271]  = 32'h3c020000;
        mem[272]  = 32'h24420138;
        mem[273]  = 32'hafc20024;
        mem[274]  = 32'h24070002;
        mem[275]  = 32'h3c020000;
        mem[276]  = 32'h24460384;
        mem[277]  = 32'h8fc40020;
        mem[278]  = 32'h8fc50024;
        mem[279]  = 32'h0c0000b2;
        mem[280]  = 32'h00000000;
        mem[281]  = 32'h00401825;
        mem[282]  = 32'h3c020000;
        mem[283]  = 32'h24420030;
        mem[284]  = 32'hac430084;
        mem[285]  = 32'h0c000076;
        mem[286]  = 32'h00000000;
        mem[287]  = 32'h00002025;
        mem[288]  = 32'h0c00005c;
        mem[289]  = 32'h00000000;
        mem[290]  = 32'h00001025;
        mem[291]  = 32'h03c0e825;
        mem[292]  = 32'h8fbf002c;
        mem[293]  = 32'h8fbe0028;
        mem[294]  = 32'h27bd0030;
        mem[295]  = 32'h03e00008;
        mem[296]  = 32'h00000000;
        mem[297]  = 32'h00000000;
        mem[298]  = 32'h00000000;
        mem[299]  = 32'h00000000;
    end
    assign data = ce ? mem[addr >> 2] : 32'b0;

endmodule
