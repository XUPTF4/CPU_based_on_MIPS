module InstMem(
        input         ce,
        input  [31:0] addr,
        output  [31:0] data
    );

    reg [31:0] mem [0:1023]; // 4KB

    initial begin
        mem[0]  = 32'h0000f025;
        mem[1]  = 32'h241d1000;
        mem[2]  = 32'h8f990028;
        mem[3]  = 32'h04110098;
        mem[4]  = 32'h00000000;
        mem[5]  = 32'h00000000;
        mem[6]  = 32'h00000000;
        mem[7]  = 32'h00000000;
        mem[8]  = 32'h10800003;
        mem[9]  = 32'h00000000;
        mem[10]  = 32'h03e00008;
        mem[11]  = 32'h00000000;
        mem[12]  = 32'h3c1c0000;
        mem[13]  = 32'h279c0000;
        mem[14]  = 32'h8f99002c;
        mem[15]  = 32'h24040001;
        mem[16]  = 32'h10000087;
        mem[17]  = 32'h00000000;
        mem[18]  = 32'h0000000c;
        mem[19]  = 32'h00000000;
        mem[20]  = 32'h03e00008;
        mem[21]  = 32'h00000000;
        mem[22]  = 32'h3c030000;
        mem[23]  = 32'h8c620040;
        mem[24]  = 32'h00000000;
        mem[25]  = 32'h24420001;
        mem[26]  = 32'h30440001;
        mem[27]  = 32'hac620040;
        mem[28]  = 32'h14800005;
        mem[29]  = 32'h00000000;
        mem[30]  = 32'h3c020000;
        mem[31]  = 32'h8c4200c8;
        mem[32]  = 32'h03e00008;
        mem[33]  = 32'h00000000;
        mem[34]  = 32'h3c020000;
        mem[35]  = 32'h8c42014c;
        mem[36]  = 32'h03e00008;
        mem[37]  = 32'h00000000;
        mem[38]  = 32'h08000016;
        mem[39]  = 32'h00000000;
        mem[40]  = 32'hafa40000;
        mem[41]  = 32'hafa50004;
        mem[42]  = 32'haca7ff8c;
        mem[43]  = 32'haca6fffc;
        mem[44]  = 32'h24a2ff7c;
        mem[45]  = 32'h03e00008;
        mem[46]  = 32'h00000000;
        mem[47]  = 32'hac040ffc;
        mem[48]  = 32'hac040ff8;
        mem[49]  = 32'h03e00008;
        mem[50]  = 32'h00000000;
        mem[51]  = 32'h27bdffe0;
        mem[52]  = 32'h3c065555;
        mem[53]  = 32'h3c02aaaa;
        mem[54]  = 32'h00801825;
        mem[55]  = 32'hafbf001c;
        mem[56]  = 32'h24050001;
        mem[57]  = 32'h24c65555;
        mem[58]  = 32'h3442aaaa;
        mem[59]  = 32'h00402025;
        mem[60]  = 32'h10650002;
        mem[61]  = 32'h00000000;
        mem[62]  = 32'h00c02025;
        mem[63]  = 32'h0c00002f;
        mem[64]  = 32'h00000000;
        mem[65]  = 32'h0c000012;
        mem[66]  = 32'h00000000;
        mem[67]  = 32'h1000fff7;
        mem[68]  = 32'h00000000;
        mem[69]  = 32'h00000000;
        mem[70]  = 32'h00000000;
        mem[71]  = 32'h00000000;
        mem[72]  = 32'h3c080000;
        mem[73]  = 32'h250300c8;
        mem[74]  = 32'h3c050000;
        mem[75]  = 32'h3c060000;
        mem[76]  = 32'h27bdffd0;
        mem[77]  = 32'h24c600cc;
        mem[78]  = 32'h00602025;
        mem[79]  = 32'h24a5014c;
        mem[80]  = 32'h24070001;
        mem[81]  = 32'hafbf002c;
        mem[82]  = 32'h0c000028;
        mem[83]  = 32'h00000000;
        mem[84]  = 32'h00a02025;
        mem[85]  = 32'h3c050000;
        mem[86]  = 32'h24070002;
        mem[87]  = 32'h24a501d0;
        mem[88]  = 32'had0200c8;
        mem[89]  = 32'h0c000028;
        mem[90]  = 32'h00000000;
        mem[91]  = 32'hac620084;
        mem[92]  = 32'h00002025;
        mem[93]  = 32'h0c000012;
        mem[94]  = 32'h00000000;
        mem[95]  = 32'h0c000008;
        mem[96]  = 32'h00000000;
        mem[97]  = 32'h8fbf002c;
        mem[98]  = 32'h00001025;
        mem[99]  = 32'h27bd0030;
        mem[100]  = 32'h03e00008;
        mem[101]  = 32'h00000000;
        mem[102]  = 32'h00000000;
        mem[103]  = 32'h00000000;
        mem[104]  = 32'h03a0d825;
        mem[105]  = 32'h27bdff7c;
        mem[106]  = 32'hafa10004;
        mem[107]  = 32'hafa20008;
        mem[108]  = 32'hafa3000c;
        mem[109]  = 32'hafa40010;
        mem[110]  = 32'hafa50014;
        mem[111]  = 32'hafa60018;
        mem[112]  = 32'hafa7001c;
        mem[113]  = 32'hafa80020;
        mem[114]  = 32'hafa90024;
        mem[115]  = 32'hafaa0028;
        mem[116]  = 32'hafab002c;
        mem[117]  = 32'hafac0030;
        mem[118]  = 32'hafad0034;
        mem[119]  = 32'hafae0038;
        mem[120]  = 32'hafaf003c;
        mem[121]  = 32'hafb00040;
        mem[122]  = 32'hafb10044;
        mem[123]  = 32'hafb20048;
        mem[124]  = 32'hafb3004c;
        mem[125]  = 32'hafb40050;
        mem[126]  = 32'hafb50054;
        mem[127]  = 32'hafb60058;
        mem[128]  = 32'hafb7005c;
        mem[129]  = 32'hafb80060;
        mem[130]  = 32'hafb90064;
        mem[131]  = 32'hafbc0070;
        mem[132]  = 32'hafbe0078;
        mem[133]  = 32'hafbf007c;
        mem[134]  = 32'hafbb0074;
        mem[135]  = 32'h03a02025;
        mem[136]  = 32'h8f990030;
        mem[137]  = 32'h0411ff9c;
        mem[138]  = 32'h00000000;
        mem[139]  = 32'h8c440010;
        mem[140]  = 32'h8c480080;
        mem[141]  = 32'h00000000;
        mem[142]  = 32'h00000000;
        mem[143]  = 32'h00000000;
        mem[144]  = 32'h00000000;
        mem[145]  = 32'h00000000;
        mem[146]  = 32'h40880000;
        mem[147]  = 32'h27bd0084;
        mem[148]  = 32'h42000018;
        mem[149]  = 32'h00000000;
        mem[150]  = 32'h00000000;
        mem[151]  = 32'h00000000;
        mem[152]  = 32'h00802025;
        mem[153]  = 32'h0000000d;
        mem[154]  = 32'h1000ffff;
        mem[155]  = 32'h00000000;
        mem[156]  = 32'h3c1c0000;
        mem[157]  = 32'h279c0000;
        mem[158]  = 32'h27bdffe0;
        mem[159]  = 32'h8f990034;
        mem[160]  = 32'hafbf001c;
        mem[161]  = 32'hafbc0010;
        mem[162]  = 32'h0411ffa5;
        mem[163]  = 32'h00000000;
        mem[164]  = 32'h00402025;
        mem[165]  = 32'h0c000098;
        mem[166]  = 32'h00000000;
        mem[167]  = 32'h00000000;
        mem[168]  = 32'h10800003;
        mem[169]  = 32'h00000000;
        mem[170]  = 32'h03e00008;
        mem[171]  = 32'h00000000;
        mem[172]  = 32'h3c1c0000;
        mem[173]  = 32'h279c0000;
        mem[174]  = 32'h8f99002c;
        mem[175]  = 32'h24040001;
        mem[176]  = 32'h1000ffe7;
        mem[177]  = 32'h00000000;
        mem[178]  = 32'h0000000c;
        mem[179]  = 32'h00000000;
        mem[180]  = 32'h03e00008;
        mem[181]  = 32'h00000000;
        mem[182]  = 32'h3c030000;
        mem[183]  = 32'h8c620040;
        mem[184]  = 32'h00000000;
        mem[185]  = 32'h24420001;
        mem[186]  = 32'h30440001;
        mem[187]  = 32'hac620040;
        mem[188]  = 32'h14800005;
        mem[189]  = 32'h00000000;
        mem[190]  = 32'h3c020000;
        mem[191]  = 32'h8c4200c8;
        mem[192]  = 32'h03e00008;
        mem[193]  = 32'h00000000;
        mem[194]  = 32'h3c020000;
        mem[195]  = 32'h8c42014c;
        mem[196]  = 32'h03e00008;
        mem[197]  = 32'h00000000;
        mem[198]  = 32'h08000016;
        mem[199]  = 32'h00000000;
        mem[200]  = 32'hafa40000;
        mem[201]  = 32'hafa50004;
        mem[202]  = 32'haca7ff8c;
        mem[203]  = 32'haca6fffc;
        mem[204]  = 32'h24a2ff7c;
        mem[205]  = 32'h03e00008;
        mem[206]  = 32'h00000000;
        mem[207]  = 32'hac040ffc;
        mem[208]  = 32'hac040ff8;
        mem[209]  = 32'h03e00008;
        mem[210]  = 32'h00000000;
        mem[211]  = 32'h27bdffe0;
        mem[212]  = 32'h3c065555;
        mem[213]  = 32'h3c02aaaa;
        mem[214]  = 32'h00801825;
        mem[215]  = 32'hafbf001c;
        mem[216]  = 32'h24050001;
        mem[217]  = 32'h24c65555;
        mem[218]  = 32'h3442aaaa;
        mem[219]  = 32'h00402025;
        mem[220]  = 32'h10650002;
        mem[221]  = 32'h00000000;
        mem[222]  = 32'h00c02025;
        mem[223]  = 32'h0c00002f;
        mem[224]  = 32'h00000000;
        mem[225]  = 32'h0c000012;
        mem[226]  = 32'h00000000;
        mem[227]  = 32'h1000fff7;
        mem[228]  = 32'h00000000;
        mem[229]  = 32'h00000000;
        mem[230]  = 32'h00000000;
        mem[231]  = 32'h00000000;
        mem[232]  = 32'h3c080000;
        mem[233]  = 32'h250300c8;
        mem[234]  = 32'h3c050000;
        mem[235]  = 32'h3c060000;
        mem[236]  = 32'h27bdffd0;
        mem[237]  = 32'h24c600cc;
        mem[238]  = 32'h00602025;
        mem[239]  = 32'h24a5014c;
        mem[240]  = 32'h24070001;
        mem[241]  = 32'hafbf002c;
        mem[242]  = 32'h0c000028;
        mem[243]  = 32'h00000000;
        mem[244]  = 32'h00a02025;
        mem[245]  = 32'h3c050000;
        mem[246]  = 32'h24070002;
        mem[247]  = 32'h24a501d0;
        mem[248]  = 32'had0200c8;
        mem[249]  = 32'h0c000028;
        mem[250]  = 32'h00000000;
        mem[251]  = 32'hac620084;
        mem[252]  = 32'h00002025;
        mem[253]  = 32'h0c000012;
        mem[254]  = 32'h00000000;
        mem[255]  = 32'h0c000008;
        mem[256]  = 32'h00000000;
        mem[257]  = 32'h8fbf002c;
        mem[258]  = 32'h00001025;
        mem[259]  = 32'h27bd0030;
        mem[260]  = 32'h03e00008;
        mem[261]  = 32'h00000000;
    end
    assign data = ce ? mem[addr >> 2] : 32'b0;

endmodule
