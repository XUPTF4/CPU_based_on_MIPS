module InstMem(
        input         ce,
        input  [31:0] addr,
        output  [31:0] data
    );

    reg [31:0] mem [0:1023]; // 4KB

    initial begin
        mem[0]  = 32'h0000f025;
        mem[1]  = 32'h241d1000;
        mem[2]  = 32'h8f990068;
        mem[3]  = 32'h041100e6;
        mem[4]  = 32'h00000000;
        mem[5]  = 32'h00000000;
        mem[6]  = 32'h00000000;
        mem[7]  = 32'h00000000;
        mem[8]  = 32'h27bdffe8;
        mem[9]  = 32'hafbe0014;
        mem[10]  = 32'h03a0f025;
        mem[11]  = 32'hafc40018;
        mem[12]  = 32'hafc5001c;
        mem[13]  = 32'hafc60020;
        mem[14]  = 32'h8fc20018;
        mem[15]  = 32'h00000000;
        mem[16]  = 32'hafc20008;
        mem[17]  = 32'h8fc2001c;
        mem[18]  = 32'h00000000;
        mem[19]  = 32'hafc2000c;
        mem[20]  = 32'h1000000c;
        mem[21]  = 32'h00000000;
        mem[22]  = 32'h8fc3000c;
        mem[23]  = 32'h00000000;
        mem[24]  = 32'h24620001;
        mem[25]  = 32'hafc2000c;
        mem[26]  = 32'h8fc20008;
        mem[27]  = 32'h00000000;
        mem[28]  = 32'h24440001;
        mem[29]  = 32'hafc40008;
        mem[30]  = 32'h80630000;
        mem[31]  = 32'h00000000;
        mem[32]  = 32'ha0430000;
        mem[33]  = 32'h8fc20020;
        mem[34]  = 32'h00000000;
        mem[35]  = 32'h2443ffff;
        mem[36]  = 32'hafc30020;
        mem[37]  = 32'h1440fff0;
        mem[38]  = 32'h00000000;
        mem[39]  = 32'h8fc20018;
        mem[40]  = 32'h03c0e825;
        mem[41]  = 32'h8fbe0014;
        mem[42]  = 32'h27bd0018;
        mem[43]  = 32'h03e00008;
        mem[44]  = 32'h00000000;
        mem[45]  = 32'h27bdffe0;
        mem[46]  = 32'hafbf001c;
        mem[47]  = 32'hafbe0018;
        mem[48]  = 32'h03a0f025;
        mem[49]  = 32'h3c1c0000;
        mem[50]  = 32'h279c0000;
        mem[51]  = 32'hafbc0010;
        mem[52]  = 32'hafc40020;
        mem[53]  = 32'h8fc20020;
        mem[54]  = 32'h00000000;
        mem[55]  = 32'h14400008;
        mem[56]  = 32'h00000000;
        mem[57]  = 32'h24040001;
        mem[58]  = 32'h8f82006c;
        mem[59]  = 32'h00000000;
        mem[60]  = 32'h0040c825;
        mem[61]  = 32'h041100a2;
        mem[62]  = 32'h00000000;
        mem[63]  = 32'h8fdc0010;
        mem[64]  = 32'h00000000;
        mem[65]  = 32'h03c0e825;
        mem[66]  = 32'h8fbf001c;
        mem[67]  = 32'h8fbe0018;
        mem[68]  = 32'h27bd0020;
        mem[69]  = 32'h03e00008;
        mem[70]  = 32'h00000000;
        mem[71]  = 32'h27bdffe8;
        mem[72]  = 32'hafbe0014;
        mem[73]  = 32'h03a0f025;
        mem[74]  = 32'hafc5001c;
        mem[75]  = 32'hafc40018;
        mem[76]  = 32'hafc70024;
        mem[77]  = 32'hafc60020;
        mem[78]  = 32'h8fc30018;
        mem[79]  = 32'h8fc20024;
        mem[80]  = 32'h00000000;
        mem[81]  = 32'h00620018;
        mem[82]  = 32'h00001012;
        mem[83]  = 32'h8fc40020;
        mem[84]  = 32'h8fc3001c;
        mem[85]  = 32'h00000000;
        mem[86]  = 32'h00830018;
        mem[87]  = 32'h00001812;
        mem[88]  = 32'h00432021;
        mem[89]  = 32'h8fc3001c;
        mem[90]  = 32'h8fc20024;
        mem[91]  = 32'h00000000;
        mem[92]  = 32'h00620019;
        mem[93]  = 32'h00001812;
        mem[94]  = 32'h00001010;
        mem[95]  = 32'h00822021;
        mem[96]  = 32'h00801025;
        mem[97]  = 32'hafc3000c;
        mem[98]  = 32'hafc20008;
        mem[99]  = 32'hafc3000c;
        mem[100]  = 32'hafc20008;
        mem[101]  = 32'h8fc3000c;
        mem[102]  = 32'h8fc20008;
        mem[103]  = 32'h03c0e825;
        mem[104]  = 32'h8fbe0014;
        mem[105]  = 32'h27bd0018;
        mem[106]  = 32'h03e00008;
        mem[107]  = 32'h00000000;
        mem[108]  = 32'h27bdffb0;
        mem[109]  = 32'hafbf004c;
        mem[110]  = 32'hafbe0048;
        mem[111]  = 32'hafb70044;
        mem[112]  = 32'hafb60040;
        mem[113]  = 32'hafb5003c;
        mem[114]  = 32'hafb40038;
        mem[115]  = 32'hafb30034;
        mem[116]  = 32'hafb20030;
        mem[117]  = 32'hafb1002c;
        mem[118]  = 32'hafb00028;
        mem[119]  = 32'h03a0f025;
        mem[120]  = 32'hafc00020;
        mem[121]  = 32'hafc00018;
        mem[122]  = 32'h10000049;
        mem[123]  = 32'h00000000;
        mem[124]  = 32'h8fc20018;
        mem[125]  = 32'h00000000;
        mem[126]  = 32'hafc2001c;
        mem[127]  = 32'h10000033;
        mem[128]  = 32'h00000000;
        mem[129]  = 32'h8fc20020;
        mem[130]  = 32'h00000000;
        mem[131]  = 32'h24430001;
        mem[132]  = 32'hafc30020;
        mem[133]  = 32'h3c040000;
        mem[134]  = 32'h000218c0;
        mem[135]  = 32'h24820010;
        mem[136]  = 32'h00621021;
        mem[137]  = 32'h8c530004;
        mem[138]  = 32'h8c520000;
        mem[139]  = 32'h3c020000;
        mem[140]  = 32'h8fc30018;
        mem[141]  = 32'h00000000;
        mem[142]  = 32'h00031880;
        mem[143]  = 32'h24420000;
        mem[144]  = 32'h00621021;
        mem[145]  = 32'h8c420000;
        mem[146]  = 32'h00000000;
        mem[147]  = 32'h0040a825;
        mem[148]  = 32'h000217c3;
        mem[149]  = 32'h0040a025;
        mem[150]  = 32'h3c020000;
        mem[151]  = 32'h8fc3001c;
        mem[152]  = 32'h00000000;
        mem[153]  = 32'h00031880;
        mem[154]  = 32'h24420000;
        mem[155]  = 32'h00621021;
        mem[156]  = 32'h8c420000;
        mem[157]  = 32'h00000000;
        mem[158]  = 32'h0040b825;
        mem[159]  = 32'h000217c3;
        mem[160]  = 32'h0040b025;
        mem[161]  = 32'h02e03825;
        mem[162]  = 32'h02c03025;
        mem[163]  = 32'h02a02825;
        mem[164]  = 32'h02802025;
        mem[165]  = 32'h0c000047;
        mem[166]  = 32'h00000000;
        mem[167]  = 32'h02428026;
        mem[168]  = 32'h02638826;
        mem[169]  = 32'h02111025;
        mem[170]  = 32'h2c420001;
        mem[171]  = 32'h304200ff;
        mem[172]  = 32'h00402025;
        mem[173]  = 32'h0c00002d;
        mem[174]  = 32'h00000000;
        mem[175]  = 32'h8fc2001c;
        mem[176]  = 32'h00000000;
        mem[177]  = 32'h24420001;
        mem[178]  = 32'hafc2001c;
        mem[179]  = 32'h8fc2001c;
        mem[180]  = 32'h00000000;
        mem[181]  = 32'h28420004;
        mem[182]  = 32'h1440ffca;
        mem[183]  = 32'h00000000;
        mem[184]  = 32'h8fc2001c;
        mem[185]  = 32'h00000000;
        mem[186]  = 32'h38420004;
        mem[187]  = 32'h2c420001;
        mem[188]  = 32'h304200ff;
        mem[189]  = 32'h00402025;
        mem[190]  = 32'h0c00002d;
        mem[191]  = 32'h00000000;
        mem[192]  = 32'h8fc20018;
        mem[193]  = 32'h00000000;
        mem[194]  = 32'h24420001;
        mem[195]  = 32'hafc20018;
        mem[196]  = 32'h8fc20018;
        mem[197]  = 32'h00000000;
        mem[198]  = 32'h28420004;
        mem[199]  = 32'h1440ffb4;
        mem[200]  = 32'h00000000;
        mem[201]  = 32'h8fc20018;
        mem[202]  = 32'h00000000;
        mem[203]  = 32'h38420004;
        mem[204]  = 32'h2c420001;
        mem[205]  = 32'h304200ff;
        mem[206]  = 32'h00402025;
        mem[207]  = 32'h0c00002d;
        mem[208]  = 32'h00000000;
        mem[209]  = 32'h00001025;
        mem[210]  = 32'h03c0e825;
        mem[211]  = 32'h8fbf004c;
        mem[212]  = 32'h8fbe0048;
        mem[213]  = 32'h8fb70044;
        mem[214]  = 32'h8fb60040;
        mem[215]  = 32'h8fb5003c;
        mem[216]  = 32'h8fb40038;
        mem[217]  = 32'h8fb30034;
        mem[218]  = 32'h8fb20030;
        mem[219]  = 32'h8fb1002c;
        mem[220]  = 32'h8fb00028;
        mem[221]  = 32'h27bd0050;
        mem[222]  = 32'h03e00008;
        mem[223]  = 32'h00000000;
        mem[224]  = 32'h27bdfff8;
        mem[225]  = 32'hafbe0004;
        mem[226]  = 32'h03a0f025;
        mem[227]  = 32'hafc40008;
        mem[228]  = 32'h8fc20008;
        mem[229]  = 32'h00000000;
        mem[230]  = 32'h00402025;
        mem[231]  = 32'h0000000d;
        mem[232]  = 32'h1000ffff;
        mem[233]  = 32'h00000000;
        mem[234]  = 32'h27bdffd8;
        mem[235]  = 32'hafbf0024;
        mem[236]  = 32'hafbe0020;
        mem[237]  = 32'h03a0f025;
        mem[238]  = 32'h3c1c0000;
        mem[239]  = 32'h279c0000;
        mem[240]  = 32'hafbc0010;
        mem[241]  = 32'h8f820070;
        mem[242]  = 32'h00000000;
        mem[243]  = 32'h0040c825;
        mem[244]  = 32'h0411ff77;
        mem[245]  = 32'h00000000;
        mem[246]  = 32'h8fdc0010;
        mem[247]  = 32'hafc20018;
        mem[248]  = 32'h8fc40018;
        mem[249]  = 32'h0c0000e0;
        mem[250]  = 32'h00000000;
        mem[251]  = 32'h8fdc0010;
        mem[252]  = 32'h00000000;
        mem[253]  = 32'h03c0e825;
        mem[254]  = 32'h8fbf0024;
        mem[255]  = 32'h8fbe0020;
        mem[256]  = 32'h27bd0028;
        mem[257]  = 32'h03e00008;
        mem[258]  = 32'h00000000;
        mem[259]  = 32'h00000000;
    end
    assign data = ce ? mem[addr >> 2] : 32'b0;

endmodule
