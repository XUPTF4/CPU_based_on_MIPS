module InstMem(
        input         ce,
        input  [31:0] addr,
        output  [31:0] data
    );

    reg [31:0] mem [0:1023]; // 4KB

    initial begin
        mem[0]  = 32'h0000f025;
        mem[1]  = 32'h241d1000;
        mem[2]  = 32'h8f990048;
        mem[3]  = 32'h04110082;
        mem[4]  = 32'h00000000;
        mem[5]  = 32'h00000000;
        mem[6]  = 32'h00000000;
        mem[7]  = 32'h00000000;
        mem[8]  = 32'h27bdffe0;
        mem[9]  = 32'hafbf001c;
        mem[10]  = 32'hafbe0018;
        mem[11]  = 32'h03a0f025;
        mem[12]  = 32'h3c1c0000;
        mem[13]  = 32'h279c0000;
        mem[14]  = 32'hafbc0010;
        mem[15]  = 32'hafc40020;
        mem[16]  = 32'h8fc20020;
        mem[17]  = 32'h00000000;
        mem[18]  = 32'h14400008;
        mem[19]  = 32'h00000000;
        mem[20]  = 32'h24040001;
        mem[21]  = 32'h8f82004c;
        mem[22]  = 32'h00000000;
        mem[23]  = 32'h0040c825;
        mem[24]  = 32'h04110063;
        mem[25]  = 32'h00000000;
        mem[26]  = 32'h8fdc0010;
        mem[27]  = 32'h00000000;
        mem[28]  = 32'h03c0e825;
        mem[29]  = 32'h8fbf001c;
        mem[30]  = 32'h8fbe0018;
        mem[31]  = 32'h27bd0020;
        mem[32]  = 32'h03e00008;
        mem[33]  = 32'h00000000;
        mem[34]  = 32'h27bdffe0;
        mem[35]  = 32'hafbf001c;
        mem[36]  = 32'hafbe0018;
        mem[37]  = 32'h03a0f025;
        mem[38]  = 32'hafc40020;
        mem[39]  = 32'h8fc20020;
        mem[40]  = 32'h00000000;
        mem[41]  = 32'h10400005;
        mem[42]  = 32'h00000000;
        mem[43]  = 32'h8fc30020;
        mem[44]  = 32'h24020001;
        mem[45]  = 32'h14620004;
        mem[46]  = 32'h00000000;
        mem[47]  = 32'h24020001;
        mem[48]  = 32'h1000000c;
        mem[49]  = 32'h00000000;
        mem[50]  = 32'h8fc20020;
        mem[51]  = 32'h00000000;
        mem[52]  = 32'h2442ffff;
        mem[53]  = 32'h00402025;
        mem[54]  = 32'h0c000022;
        mem[55]  = 32'h00000000;
        mem[56]  = 32'h00401825;
        mem[57]  = 32'h8fc20020;
        mem[58]  = 32'h00000000;
        mem[59]  = 32'h00620018;
        mem[60]  = 32'h00001012;
        mem[61]  = 32'h03c0e825;
        mem[62]  = 32'h8fbf001c;
        mem[63]  = 32'h8fbe0018;
        mem[64]  = 32'h27bd0020;
        mem[65]  = 32'h03e00008;
        mem[66]  = 32'h00000000;
        mem[67]  = 32'h27bdffd8;
        mem[68]  = 32'hafbf0024;
        mem[69]  = 32'hafbe0020;
        mem[70]  = 32'h03a0f025;
        mem[71]  = 32'hafc00018;
        mem[72]  = 32'h10000025;
        mem[73]  = 32'h00000000;
        mem[74]  = 32'h8fc40018;
        mem[75]  = 32'h0c000022;
        mem[76]  = 32'h00000000;
        mem[77]  = 32'h00402025;
        mem[78]  = 32'h3c020000;
        mem[79]  = 32'h8fc30018;
        mem[80]  = 32'h00000000;
        mem[81]  = 32'h00031880;
        mem[82]  = 32'h24420060;
        mem[83]  = 32'h00621021;
        mem[84]  = 32'hac440000;
        mem[85]  = 32'h3c020000;
        mem[86]  = 32'h8fc30018;
        mem[87]  = 32'h00000000;
        mem[88]  = 32'h00031880;
        mem[89]  = 32'h24420060;
        mem[90]  = 32'h00621021;
        mem[91]  = 32'h8c430000;
        mem[92]  = 32'h3c020000;
        mem[93]  = 32'h8fc40018;
        mem[94]  = 32'h00000000;
        mem[95]  = 32'h00042080;
        mem[96]  = 32'h24420000;
        mem[97]  = 32'h00821021;
        mem[98]  = 32'h8c420000;
        mem[99]  = 32'h00000000;
        mem[100]  = 32'h00621026;
        mem[101]  = 32'h2c420001;
        mem[102]  = 32'h304200ff;
        mem[103]  = 32'h00402025;
        mem[104]  = 32'h0c000008;
        mem[105]  = 32'h00000000;
        mem[106]  = 32'h8fc20018;
        mem[107]  = 32'h00000000;
        mem[108]  = 32'h24420001;
        mem[109]  = 32'hafc20018;
        mem[110]  = 32'h8fc20018;
        mem[111]  = 32'h00000000;
        mem[112]  = 32'h2842000d;
        mem[113]  = 32'h1440ffd8;
        mem[114]  = 32'h00000000;
        mem[115]  = 32'h00001025;
        mem[116]  = 32'h03c0e825;
        mem[117]  = 32'h8fbf0024;
        mem[118]  = 32'h8fbe0020;
        mem[119]  = 32'h27bd0028;
        mem[120]  = 32'h03e00008;
        mem[121]  = 32'h00000000;
        mem[122]  = 32'h00000000;
        mem[123]  = 32'h00000000;
        mem[124]  = 32'h27bdfff8;
        mem[125]  = 32'hafbe0004;
        mem[126]  = 32'h03a0f025;
        mem[127]  = 32'hafc40008;
        mem[128]  = 32'h8fc20008;
        mem[129]  = 32'h00000000;
        mem[130]  = 32'h00402025;
        mem[131]  = 32'h0000000d;
        mem[132]  = 32'h1000ffff;
        mem[133]  = 32'h00000000;
        mem[134]  = 32'h27bdffd8;
        mem[135]  = 32'hafbf0024;
        mem[136]  = 32'hafbe0020;
        mem[137]  = 32'h03a0f025;
        mem[138]  = 32'h3c1c0000;
        mem[139]  = 32'h279c0000;
        mem[140]  = 32'hafbc0010;
        mem[141]  = 32'h8f820050;
        mem[142]  = 32'h00000000;
        mem[143]  = 32'h0040c825;
        mem[144]  = 32'h0411ffb2;
        mem[145]  = 32'h00000000;
        mem[146]  = 32'h8fdc0010;
        mem[147]  = 32'hafc20018;
        mem[148]  = 32'h8fc40018;
        mem[149]  = 32'h0c00007c;
        mem[150]  = 32'h00000000;
        mem[151]  = 32'h8fdc0010;
        mem[152]  = 32'h00000000;
        mem[153]  = 32'h03c0e825;
        mem[154]  = 32'h8fbf0024;
        mem[155]  = 32'h8fbe0020;
        mem[156]  = 32'h27bd0028;
        mem[157]  = 32'h03e00008;
        mem[158]  = 32'h00000000;
        mem[159]  = 32'h00000000;
    end
    assign data = ce ? mem[addr >> 2] : 32'b0;

endmodule
