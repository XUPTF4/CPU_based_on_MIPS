// 运算单元
// 这里主要实现 ALU
// 发出跳转信号：跳转信号的生成需要 ALU，放在 IDU 是不合理的

`include "Helpers.v"  // 包含 constants.v 文件
module EXU (
        input wire [31:0] regaData_i,         // 源 A 数据
        input wire [31:0] regbData_i,         // 源 B 数据
        // input wire  regcWr_i,               // 写使能
        // input wire [4:0] regcAddr_i,        // 寄存器写地址

        // for reg
        output reg [31:0] regcData,         // 寄存器写数据
        output wire [4:0] regcAddr,         // 寄存器写地址
        output wire regcWr,                   // 寄存器写使能
        output wire [1:0] WB_SEL,      // WB 数据来源 (输入信号)
        output wire [0:0] REG_EN,      // 寄存器写使能 (输入信号)

        output reg [31:0] jAddr, 	        // 跳转地址

        // for mem
        output wire [31:0] memAddr,         // 内存访问地址
        output wire [31:0] memData,         // 内存写数据
        output wire readWr,                 // 内存读使能
        output wire writeWr,                // 内存写使能
        output wire [3:0] rmask,            // 读掩码
        output wire [3:0] wmask,            // 写掩码


        // 来自上游的信号
        input wire [5:0] EXE_FUNC_i,    // ALU 功能 (输入信号)
        input wire [0:0] W_MEM_EN_i,      // 内存写使能 (输入信号)
        input wire [0:0] R_MEM_EN_i,      // 内存读使能 (输入信号)
        input wire [3:0] W_MASK_i,      // w_mask (输入信号)
        input wire [3:0] R_MASK_i,      // r_mask (输入信号)
        input wire [0:0] REG_EN_i,      // 寄存器写使能 (输入信号)
        input wire [1:0] WB_SEL_i,      // WB 数据来源 (输入信号)
        input wire [4:0] Reg_Target_i,     // WB 数据地址
        input wire [31:0] rt_data_o     // store 指令写入的数据，for MEM
    );

    // WB
    assign regcData = alu_out;
    assign regcAddr = Reg_Target_i;
    assign regcWr = R_MEM_EN_i;
    assign REG_EN = REG_EN_i;
    assign WB_SEL = WB_SEL_i;

    // 跳转地址
    assign jAddr = 32'd0;

    // 内存信号
    assign memAddr = alu_out; // 如果是 load：OK；如果是 store：
    assign memData = rt_data_o; // 那也 OK
    assign readWr = R_MEM_EN_i;
    assign writeWr = W_MEM_EN_i;
    assign rmask = R_MASK_i;
    assign wmask = W_MASK_i;


    reg [31:0] alu_out;
    // ALU
    always @(*) begin
        case (EXE_FUNC_i)
            ALU_ADD:
                alu_out = regaData_i + regbData_i;
            ALU_LW:
                alu_out = regaData_i + regbData_i; // LW
            ALU_SW:
                alu_out = regaData_i + regbData_i; // SW
            ALU_JAL:
                alu_out = regaData_i + regbData_i; // JAL
            ALU_BEQ:
                alu_out = (regaData_i << 2) + regbData_i;
            ALU_BNE:
                alu_out = (regaData_i << 2) + regbData_i;
            ALU_SUB:
                alu_out = regaData_i - regbData_i;
            ALU_AND:
                alu_out = regaData_i & regbData_i;
            ALU_OR:
                alu_out = regaData_i | regbData_i;
            ALU_XOR:
                alu_out = regaData_i ^ regbData_i;
            ALU_SLL:
                alu_out = regbData_i << regaData_i;
            ALU_SRL:
                alu_out = regbData_i >> regaData_i;
            ALU_SRA:
                alu_out = regbData_i >>> regaData_i; // 数学右移
            ALU_LUI:
                alu_out = regaData_i;
            default:
                alu_out = 32'b0;
        endcase
    end


    always @(*) begin
        case (EXE_FUNC_i)
            ALU_J:
                jAddr = {regaData_i[31:28],regbData_i[25:0],2'b00};
            ALU_JR:
                jAddr = {regaData_i[31:28],regbData_i[25:0],2'b00};
            ALU_JAL:
                jAddr = {regaData_i[31:28],regbData_i[25:0],2'b00};
            ALU_BEQ:
                jAddr = alu_out; // 直接连接 alu_out
            ALU_BNE:
                jAddr = alu_out; // 直接连接 alu_out
            default:
                jAddr = 32'b0;
        endcase
    end
endmodule
