module InstMem(
        input         ce,
        input  [31:0] addr,
        output  [31:0] data
    );

    reg [31:0] mem [0:1023]; // 4KB

    initial begin
        mem[0]  = 32'h0000f025;
        mem[1]  = 32'h241d1000;
        mem[2]  = 32'h8f990028;
        mem[3]  = 32'h04110088;
        mem[4]  = 32'h00000000;
        mem[5]  = 32'h00000000;
        mem[6]  = 32'h00000000;
        mem[7]  = 32'h00000000;
        mem[8]  = 32'h10800003;
        mem[9]  = 32'h00000000;
        mem[10]  = 32'h03e00008;
        mem[11]  = 32'h00000000;
        mem[12]  = 32'h3c1c0000;
        mem[13]  = 32'h24040001;
        mem[14]  = 32'h279c0000;
        mem[15]  = 32'h8f99002c;
        mem[16]  = 32'h10000077;
        mem[17]  = 32'h00000000;
        mem[18]  = 32'h0000000c;
        mem[19]  = 32'h00000000;
        mem[20]  = 32'h03e00008;
        mem[21]  = 32'h00000000;
        mem[22]  = 32'h3c020000;
        mem[23]  = 32'h8c420000;
        mem[24]  = 32'h8c420000;
        mem[25]  = 32'hac400000;
        mem[26]  = 32'hac410004;
        mem[27]  = 32'hac420008;
        mem[28]  = 32'hac43000c;
        mem[29]  = 32'hac440010;
        mem[30]  = 32'h03e00008;
        mem[31]  = 32'h00000000;
        mem[32]  = 32'h3c020000;
        mem[33]  = 32'h8c430000;
        mem[34]  = 32'h8c630000;
        mem[35]  = 32'h8c600000;
        mem[36]  = 32'h8c610004;
        mem[37]  = 32'h8c620008;
        mem[38]  = 32'h8c63000c;
        mem[39]  = 32'h8c640010;
        mem[40]  = 32'h8c420000;
        mem[41]  = 32'h8c420000;
        mem[42]  = 32'h8c480080;
        mem[43]  = 32'h40887000;
        mem[44]  = 32'h03e00008;
        mem[45]  = 32'h00000000;
        mem[46]  = 32'h3c030000;
        mem[47]  = 32'h3c020000;
        mem[48]  = 32'h8c640000;
        mem[49]  = 32'h244200c4;
        mem[50]  = 32'h10820004;
        mem[51]  = 32'h00000000;
        mem[52]  = 32'hac620000;
        mem[53]  = 32'h03e00008;
        mem[54]  = 32'h00000000;
        mem[55]  = 32'h3c020000;
        mem[56]  = 32'h24420148;
        mem[57]  = 32'hac620000;
        mem[58]  = 32'h03e00008;
        mem[59]  = 32'h00000000;
        mem[60]  = 32'h27bdffe0;
        mem[61]  = 32'hafbf001c;
        mem[62]  = 32'h0c000016;
        mem[63]  = 32'h00000000;
        mem[64]  = 32'h0c00002e;
        mem[65]  = 32'h00000000;
        mem[66]  = 32'h0c000020;
        mem[67]  = 32'h00000000;
        mem[68]  = 32'h42000018;
        mem[69]  = 32'h8fbf001c;
        mem[70]  = 32'h27bd0020;
        mem[71]  = 32'h03e00008;
        mem[72]  = 32'h00000000;
        mem[73]  = 32'h24a2ff7c;
        mem[74]  = 32'hafa40000;
        mem[75]  = 32'hafa50004;
        mem[76]  = 32'haca6fffc;
        mem[77]  = 32'haca7ff8c;
        mem[78]  = 32'h03e00008;
        mem[79]  = 32'h00000000;
        mem[80]  = 32'hac040ffc;
        mem[81]  = 32'h03e00008;
        mem[82]  = 32'h00000000;
        mem[83]  = 32'h27bdffe0;
        mem[84]  = 32'h3c07bbbb;
        mem[85]  = 32'h3c03aaaa;
        mem[86]  = 32'h24060001;
        mem[87]  = 32'hafbf001c;
        mem[88]  = 32'h00802825;
        mem[89]  = 32'h34e7bbbb;
        mem[90]  = 32'h3463aaaa;
        mem[91]  = 32'h8ca20000;
        mem[92]  = 32'h00602025;
        mem[93]  = 32'h10460002;
        mem[94]  = 32'h00000000;
        mem[95]  = 32'h00e02025;
        mem[96]  = 32'h0c000050;
        mem[97]  = 32'h00000000;
        mem[98]  = 32'h0c000012;
        mem[99]  = 32'h00000000;
        mem[100]  = 32'h1000fff6;
        mem[101]  = 32'h00000000;
        mem[102]  = 32'h00000000;
        mem[103]  = 32'h00000000;
        mem[104]  = 32'h3c090000;
        mem[105]  = 32'h3c030000;
        mem[106]  = 32'h3c060000;
        mem[107]  = 32'h27bdffd0;
        mem[108]  = 32'h24630148;
        mem[109]  = 32'h252800c4;
        mem[110]  = 32'h24c6014c;
        mem[111]  = 32'hafbf002c;
        mem[112]  = 32'h24070001;
        mem[113]  = 32'h01002025;
        mem[114]  = 32'h00602825;
        mem[115]  = 32'h0c000049;
        mem[116]  = 32'h00000000;
        mem[117]  = 32'h3c050000;
        mem[118]  = 32'h24070002;
        mem[119]  = 32'had2200c4;
        mem[120]  = 32'h24a501cc;
        mem[121]  = 32'h00602025;
        mem[122]  = 32'h0c000049;
        mem[123]  = 32'h00000000;
        mem[124]  = 32'h00002025;
        mem[125]  = 32'had020084;
        mem[126]  = 32'h0c000012;
        mem[127]  = 32'h00000000;
        mem[128]  = 32'h0c000008;
        mem[129]  = 32'h00000000;
        mem[130]  = 32'h00001025;
        mem[131]  = 32'h8fbf002c;
        mem[132]  = 32'h27bd0030;
        mem[133]  = 32'h03e00008;
        mem[134]  = 32'h00000000;
        mem[135]  = 32'h00000000;
        mem[136]  = 32'h00802025;
        mem[137]  = 32'h0000000d;
        mem[138]  = 32'h1000ffff;
        mem[139]  = 32'h00000000;
        mem[140]  = 32'h3c1c0000;
        mem[141]  = 32'h27bdffe0;
        mem[142]  = 32'h279c0000;
        mem[143]  = 32'hafbf001c;
        mem[144]  = 32'hafbc0010;
        mem[145]  = 32'h8f990030;
        mem[146]  = 32'h0411ffd5;
        mem[147]  = 32'h00000000;
        mem[148]  = 32'h00402025;
        mem[149]  = 32'h0c000088;
        mem[150]  = 32'h00000000;
        mem[151]  = 32'h00000000;
        mem[152]  = 32'h10800003;
        mem[153]  = 32'h00000000;
        mem[154]  = 32'h03e00008;
        mem[155]  = 32'h00000000;
        mem[156]  = 32'h3c1c0000;
        mem[157]  = 32'h24040001;
        mem[158]  = 32'h279c0000;
        mem[159]  = 32'h8f99002c;
        mem[160]  = 32'h1000ffe7;
        mem[161]  = 32'h00000000;
        mem[162]  = 32'h0000000c;
        mem[163]  = 32'h00000000;
        mem[164]  = 32'h03e00008;
        mem[165]  = 32'h00000000;
        mem[166]  = 32'h3c020000;
        mem[167]  = 32'h8c420000;
        mem[168]  = 32'h8c420000;
        mem[169]  = 32'hac400000;
        mem[170]  = 32'hac410004;
        mem[171]  = 32'hac420008;
        mem[172]  = 32'hac43000c;
        mem[173]  = 32'hac440010;
        mem[174]  = 32'h03e00008;
        mem[175]  = 32'h00000000;
        mem[176]  = 32'h3c020000;
        mem[177]  = 32'h8c430000;
        mem[178]  = 32'h8c630000;
        mem[179]  = 32'h8c600000;
        mem[180]  = 32'h8c610004;
        mem[181]  = 32'h8c620008;
        mem[182]  = 32'h8c63000c;
        mem[183]  = 32'h8c640010;
        mem[184]  = 32'h8c420000;
        mem[185]  = 32'h8c420000;
        mem[186]  = 32'h8c480080;
        mem[187]  = 32'h40887000;
        mem[188]  = 32'h03e00008;
        mem[189]  = 32'h00000000;
        mem[190]  = 32'h3c030000;
        mem[191]  = 32'h3c020000;
        mem[192]  = 32'h8c640000;
        mem[193]  = 32'h244200c4;
        mem[194]  = 32'h10820004;
        mem[195]  = 32'h00000000;
        mem[196]  = 32'hac620000;
        mem[197]  = 32'h03e00008;
        mem[198]  = 32'h00000000;
        mem[199]  = 32'h3c020000;
        mem[200]  = 32'h24420148;
        mem[201]  = 32'hac620000;
        mem[202]  = 32'h03e00008;
        mem[203]  = 32'h00000000;
        mem[204]  = 32'h27bdffe0;
        mem[205]  = 32'hafbf001c;
        mem[206]  = 32'h0c000016;
        mem[207]  = 32'h00000000;
        mem[208]  = 32'h0c00002e;
        mem[209]  = 32'h00000000;
        mem[210]  = 32'h0c000020;
        mem[211]  = 32'h00000000;
        mem[212]  = 32'h42000018;
        mem[213]  = 32'h8fbf001c;
        mem[214]  = 32'h27bd0020;
        mem[215]  = 32'h03e00008;
        mem[216]  = 32'h00000000;
        mem[217]  = 32'h24a2ff7c;
        mem[218]  = 32'hafa40000;
        mem[219]  = 32'hafa50004;
        mem[220]  = 32'haca6fffc;
        mem[221]  = 32'haca7ff8c;
        mem[222]  = 32'h03e00008;
        mem[223]  = 32'h00000000;
        mem[224]  = 32'hac040ffc;
        mem[225]  = 32'h03e00008;
        mem[226]  = 32'h00000000;
        mem[227]  = 32'h27bdffe0;
        mem[228]  = 32'h3c07bbbb;
        mem[229]  = 32'h3c03aaaa;
        mem[230]  = 32'h24060001;
        mem[231]  = 32'hafbf001c;
        mem[232]  = 32'h00802825;
        mem[233]  = 32'h34e7bbbb;
        mem[234]  = 32'h3463aaaa;
        mem[235]  = 32'h8ca20000;
        mem[236]  = 32'h00602025;
        mem[237]  = 32'h10460002;
        mem[238]  = 32'h00000000;
        mem[239]  = 32'h00e02025;
        mem[240]  = 32'h0c000050;
        mem[241]  = 32'h00000000;
        mem[242]  = 32'h0c000012;
        mem[243]  = 32'h00000000;
        mem[244]  = 32'h1000fff6;
        mem[245]  = 32'h00000000;
        mem[246]  = 32'h00000000;
        mem[247]  = 32'h00000000;
        mem[248]  = 32'h3c090000;
        mem[249]  = 32'h3c030000;
        mem[250]  = 32'h3c060000;
        mem[251]  = 32'h27bdffd0;
        mem[252]  = 32'h24630148;
        mem[253]  = 32'h252800c4;
        mem[254]  = 32'h24c6014c;
        mem[255]  = 32'hafbf002c;
        mem[256]  = 32'h24070001;
        mem[257]  = 32'h01002025;
        mem[258]  = 32'h00602825;
        mem[259]  = 32'h0c000049;
        mem[260]  = 32'h00000000;
        mem[261]  = 32'h3c050000;
        mem[262]  = 32'h24070002;
        mem[263]  = 32'had2200c4;
        mem[264]  = 32'h24a501cc;
        mem[265]  = 32'h00602025;
        mem[266]  = 32'h0c000049;
        mem[267]  = 32'h00000000;
        mem[268]  = 32'h00002025;
        mem[269]  = 32'had020084;
        mem[270]  = 32'h0c000012;
        mem[271]  = 32'h00000000;
        mem[272]  = 32'h0c000008;
        mem[273]  = 32'h00000000;
        mem[274]  = 32'h00001025;
        mem[275]  = 32'h8fbf002c;
        mem[276]  = 32'h27bd0030;
        mem[277]  = 32'h03e00008;
        mem[278]  = 32'h00000000;
    end
    assign data = ce ? mem[addr >> 2] : 32'b0;

endmodule
